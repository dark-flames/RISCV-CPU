`define LITTLE_ENDIAN	1
//`define ST_DEBUG	1
//`define LD_DEBUG	1
//`define VCD		1
